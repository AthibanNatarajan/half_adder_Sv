interface haif();
logic a;
logic b;
logic sum;
logic cout;
endinterface
